module mkTest ();

  rule hello;
    $display("Hello");
    $finish();
  endrule

endmodule
